module tx (
    input clk,
    input rst,
    input tx_ready,
    input [7:0] tx_data,
    output reg tx,
    output reg tx_rd
);
  parameter DIV_CNT = 10'd867;
  parameter HDIV_CNT = 10'd433;
  parameter TX_CNT = 4'h9;
  parameter C_IDLE = 1'b0;
  parameter C_TX = 1'b1;
  reg curr_state, next_state;
  reg [9:0] div_cnt;
  reg [4:0] tx_cnt;
  reg [7:0] tx_reg;

  initial begin
    curr_state = C_IDLE;
    div_cnt = 10'h0;
    tx_cnt = 4'h0;
    tx_rd = 1'b0;
    tx_reg = 8'h0;
    tx = 1'b1;
  end

  always @(posedge clk or posedge rst) begin
    if (rst) curr_state <= C_IDLE;
    else curr_state <= next_state;
  end
  always @(*) begin
    case (curr_state)
      C_IDLE:
      if (tx_ready == 1'b1) next_state = C_TX;
      else next_state = C_IDLE;
      C_TX:
      if ((div_cnt == DIV_CNT) && (tx_cnt >= TX_CNT)) next_state = C_IDLE;
      else next_state = C_TX;
    endcase
  end
  always @(posedge clk or posedge rst) begin
    if (rst) div_cnt <= 10'h0;
    else if (curr_state == C_TX) begin
      if (div_cnt >= DIV_CNT) div_cnt <= 10'h0;
      else div_cnt <= div_cnt + 10'h1;
    end else div_cnt <= 10'h0;
  end
  always @(posedge clk or posedge rst) begin
    if (rst) tx_cnt <= 4'h0;
    else if (curr_state == C_TX) begin
      if (div_cnt == DIV_CNT) tx_cnt <= tx_cnt + 1'b1;
    end else tx_cnt <= 4'h0;
  end
  always @(posedge clk or posedge rst) begin
    if (rst) tx_rd <= 1'b0;
    else if ((curr_state == C_IDLE) && (tx_ready == 1'b1)) tx_rd <= 1'b1;
    else tx_rd <= 1'b0;
  end
  always @(posedge clk or posedge rst) begin
    if (rst) tx_reg <= 8'b0;
    else if ((curr_state == C_IDLE) && (tx_ready == 1'b1)) tx_reg <= tx_data;
  end
  always @(posedge clk or posedge rst) begin
    if (rst) tx <= 1'b1;
    else if (curr_state == C_IDLE) tx <= 1'b1;
    else if (div_cnt == 10'h0) begin
      case (tx_cnt)
        4'h0: tx <= 1'b0;
        4'h1: tx <= tx_reg[0];
        4'h2: tx <= tx_reg[1];
        4'h3: tx <= tx_reg[2];
        4'h4: tx <= tx_reg[3];
        4'h5: tx <= tx_reg[4];
        4'h6: tx <= tx_reg[5];
        4'h7: tx <= tx_reg[6];
        4'h8: tx <= tx_reg[7];
        4'h9: tx <= 1'b1;
      endcase
    end
  end
endmodule